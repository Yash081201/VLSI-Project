NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

DIVIDERCHAR "/" ;

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.042 ;
  SPACING 0.09 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M1

LAYER V1
  TYPE CUT ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M2

LAYER V2
  TYPE CUT ;
END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M3

LAYER V3
  TYPE CUT ;
END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M4

LAYER V4
  TYPE CUT ;
END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
END M5

LAYER V5
  TYPE CUT ;
END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.26 0.26 ;
  WIDTH 0.14 ;
  AREA 0.052 ;
  SPACING 0.1 ;
  SPACING 0.19 RANGE 1.76 4 ;
  SPACING 0.29 RANGE 4 8 ;
  SPACING 1.05 RANGE 8 25 ;
  SPACING 1.85 RANGE 25 100000 ;
  END M6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

SPACING
  SAMENET M1  M1    0.09 STACK ;
  SAMENET M2  M2    0.1 STACK ;
  SAMENET M3  M3    0.1 STACK ;
  SAMENET M4  M4    0.1 STACK ;
  SAMENET M5  M5    0.1 STACK ;
  SAMENET M6  M6    0.1 STACK ;
  SAMENET V1  V1    0.1 ;
  SAMENET V2  V2    0.1 ;
  SAMENET V3  V3    0.1 ;
  SAMENET V4  V4    0.1 ;
  SAMENET V5  V5    0.1 ;
  SAMENET V1  V2    0.00 STACK ;
  SAMENET V2  V3    0.00 STACK ;
  SAMENET V3  V4    0.00 STACK ;
  SAMENET V4  V5    0.00 STACK ;
  SAMENET V1  V3    0.00 STACK ;
  SAMENET V2  V4    0.00 STACK ;
  SAMENET V3  V5    0.00 STACK ;
  SAMENET V1  V4    0.00 STACK ;
  SAMENET V2  V5    0.00 STACK ;
  SAMENET V1  V5    0.00 STACK ;
END SPACING


VIA via5 DEFAULT
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via5

VIA via4 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via4

VIA via3 DEFAULT
  LAYER M4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via3

VIA via2 DEFAULT
  LAYER M3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via2

VIA via1 DEFAULT
  LAYER M2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
END via1


VIARULE via1Array GENERATE
  LAYER M1 ;
  DIRECTION HORIZONTAL ;
  OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via1Array


VIARULE via2Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M2 ;
  DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via2Array


VIARULE via3Array GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via3Array

VIARULE via4Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER V4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via4Array

VIARULE via5Array GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
    OVERHANG 0.03 ;
    METALOVERHANG 0 ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
    OVERHANG 0.045 ;
    METALOVERHANG 0 ;
  LAYER V5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END via5Array

VIARULE TURNM1 GENERATE
  LAYER M1 ;
    DIRECTION HORIZONTAL ;
  LAYER M1 ;
    DIRECTION VERTICAL ;
END TURNM1

VIARULE TURNM2 GENERATE
  LAYER M2 ;
    DIRECTION HORIZONTAL ;
  LAYER M2 ;
    DIRECTION VERTICAL ;
END TURNM2

VIARULE TURNM3 GENERATE
  LAYER M3 ;
    DIRECTION HORIZONTAL ;
  LAYER M3 ;
    DIRECTION VERTICAL ;
END TURNM3

VIARULE TURNM4 GENERATE
  LAYER M4 ;
    DIRECTION HORIZONTAL ;
  LAYER M4 ;
    DIRECTION VERTICAL ;
END TURNM4

VIARULE TURNM5 GENERATE
  LAYER M5 ;
    DIRECTION HORIZONTAL ;
  LAYER M5 ;
    DIRECTION VERTICAL ;
END TURNM5

VIARULE TURNM6 GENERATE
  LAYER M6 ;
    DIRECTION HORIZONTAL ;
  LAYER M6 ;
    DIRECTION VERTICAL ;
END TURNM6


SITE  CoreSite
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.9 ;
END  CoreSite

SITE  TDCoverSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  TDCoverSite

SITE  SBlockSite
    CLASS       CORE ;
    SIZE        0.0500 BY 0.0500 ;
END  SBlockSite

SITE  PortCellSite
    CLASS       PAD ;
    SIZE        0.0500 BY 0.0500 ;
END  PortCellSite

SITE  Core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SYMMETRY    X ;
    SIZE        0.260 BY 4.9 ;
END  Core


MACRO AOI21
  CLASS CORE ;
  ORIGIN -7.636 -4.63 ;
  FOREIGN AOI21 7.636 4.63 ;
  SIZE 2.64 BY 5.06 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.761 6.878 8.871 7.261 ;
      LAYER M2 ;
        RECT 8.741 6.872 8.871 7.272 ;
      LAYER V1 ;
        RECT 8.766 7.024 8.866 7.124 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 8.161 6.878 8.271 7.261 ;
      LAYER M2 ;
        RECT 8.141 6.872 8.271 7.272 ;
      LAYER V1 ;
        RECT 8.166 7.024 8.266 7.124 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.361 6.878 9.471 7.261 ;
      LAYER M2 ;
        RECT 9.341 6.872 9.471 7.272 ;
      LAYER V1 ;
        RECT 9.366 7.024 9.466 7.124 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.64 6.866 9.756 7.264 ;
        RECT 9.64 6.654 9.73 8.331 ;
        RECT 9.081 6.654 9.73 6.744 ;
        RECT 9.081 5.964 9.171 6.744 ;
      LAYER M2 ;
        RECT 9.641 6.878 9.771 7.278 ;
      LAYER V1 ;
        RECT 9.645 7.033 9.745 7.133 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 7.756 9.41 10.156 9.53 ;
        RECT 8.391 7.531 8.481 9.53 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 7.756 4.63 10.156 4.75 ;
        RECT 9.495 4.63 9.585 6.564 ;
        RECT 8.126 4.63 8.216 6.564 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 9.081 7.351 9.171 8.331 ;
      RECT 8.126 7.351 8.216 8.331 ;
      RECT 8.126 7.351 9.171 7.441 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END AOI21

MACRO AOI22
  CLASS CORE ;
  ORIGIN -9.721 -5.653 ;
  FOREIGN AOI22 9.721 5.653 ;
  SIZE 2.7 BY 4.901 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.706 7.865 10.821 8.265 ;
      LAYER M2 ;
        RECT 10.706 7.895 10.836 8.295 ;
      LAYER V1 ;
        RECT 10.715 8.05 10.815 8.15 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.121 7.865 10.236 8.265 ;
      LAYER M2 ;
        RECT 10.106 7.895 10.236 8.295 ;
      LAYER V1 ;
        RECT 10.126 8.05 10.226 8.15 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.306 7.865 11.421 8.265 ;
      LAYER M2 ;
        RECT 11.306 7.895 11.436 8.295 ;
      LAYER V1 ;
        RECT 11.315 8.05 11.415 8.15 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.906 7.865 12.021 8.265 ;
      LAYER M2 ;
        RECT 11.906 7.895 12.036 8.295 ;
      LAYER V1 ;
        RECT 11.915 8.05 12.015 8.15 ;
    END
  END D
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.406 7.658 11.009 7.755 ;
        RECT 10.919 6.987 11.009 7.755 ;
        RECT 10.406 7.865 10.521 8.265 ;
        RECT 10.406 7.658 10.496 9.354 ;
      LAYER M2 ;
        RECT 10.406 7.894 10.536 8.294 ;
      LAYER V1 ;
        RECT 10.416 8.049 10.516 8.149 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 9.721 10.433 12.421 10.553 ;
        RECT 11.426 8.554 11.516 10.553 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 9.721 5.653 12.421 5.773 ;
        RECT 12.026 5.653 12.116 7.587 ;
        RECT 10.091 5.653 10.181 7.587 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 10.091 9.594 10.949 9.684 ;
      RECT 10.859 8.374 10.949 9.684 ;
      RECT 10.091 8.554 10.181 9.684 ;
      RECT 12.026 8.374 12.116 9.354 ;
      RECT 10.859 8.374 12.116 8.464 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END AOI22

MACRO DFF
  CLASS CORE ;
  ORIGIN -8.44 -7.139 ;
  FOREIGN DFF 8.44 7.139 ;
  SIZE 5.1 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 13.045 9.351 13.155 9.751 ;
      LAYER M2 ;
        RECT 13.025 9.381 13.155 9.781 ;
      LAYER V1 ;
        RECT 13.05 9.533 13.15 9.633 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.045 9.351 10.155 9.751 ;
      LAYER M2 ;
        RECT 10.025 9.381 10.155 9.781 ;
      LAYER V1 ;
        RECT 10.05 9.533 10.15 9.633 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.443 9.351 12.555 9.751 ;
        RECT 12.443 8.473 12.533 10.84 ;
      LAYER M2 ;
        RECT 12.425 9.381 12.555 9.781 ;
      LAYER V1 ;
        RECT 12.45 9.533 12.55 9.633 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.44 11.919 13.54 12.039 ;
        RECT 12.875 10.04 12.965 12.039 ;
        RECT 11.76 10.04 11.85 12.039 ;
        RECT 10.185 10.04 10.275 12.039 ;
        RECT 8.925 10.04 9.015 12.039 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.44 7.139 13.54 7.259 ;
        RECT 12.875 7.139 12.965 9.073 ;
        RECT 11.76 7.139 11.85 9.073 ;
        RECT 10.196 7.139 10.286 9.073 ;
        RECT 8.925 7.139 9.015 9.073 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 13.245 11.328 13.4 11.486 ;
      RECT 13.305 8.473 13.395 11.486 ;
      RECT 12.09 11.095 12.245 11.253 ;
      RECT 12.12 8.058 12.21 11.253 ;
      RECT 12.09 8.058 12.24 8.208 ;
      RECT 11.08 8.473 11.17 10.84 ;
      RECT 11.862 9.657 12.011 9.806 ;
      RECT 11.08 9.687 12.011 9.777 ;
      RECT 11.178 11.098 11.362 11.258 ;
      RECT 9.61 11.113 9.95 11.243 ;
      RECT 9.86 8.201 9.95 11.243 ;
      RECT 10.668 11.133 11.362 11.223 ;
      RECT 10.668 9.145 10.759 11.223 ;
      RECT 9.762 9.163 10.759 9.253 ;
      RECT 9.331 8.167 9.492 8.325 ;
      RECT 9.331 8.201 9.95 8.291 ;
      RECT 9.497 8.473 9.587 10.84 ;
      RECT 8.774 9.653 8.919 9.812 ;
      RECT 8.774 9.687 9.587 9.777 ;
      RECT 8.585 7.788 8.675 10.84 ;
      RECT 8.55 7.788 8.726 7.983 ;
  END
END DFF

MACRO Filler_ckt
  CLASS CORE ;
  ORIGIN -7.804 -5.758 ;
  FOREIGN Filler_ckt 7.804 5.758 ;
  SIZE 0.3 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 7.779 10.538 8.129 10.658 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 7.779 5.758 8.129 5.878 ;
    END
  END VSS
  PROPERTY CatenaDesignType "deviceLevel" ;
END Filler_ckt

MACRO INVERTER
  CLASS CORE ;
  ORIGIN -11.643 -5.787 ;
  FOREIGN INVERTER 11.643 5.787 ;
  SIZE 1.2 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.048 8.008 12.158 8.393 ;
      LAYER M2 ;
        RECT 12.028 8.029 12.158 8.429 ;
      LAYER V1 ;
        RECT 12.049 8.174 12.149 8.274 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.328 7.999 12.443 8.399 ;
        RECT 12.328 7.121 12.418 9.488 ;
      LAYER M2 ;
        RECT 12.328 8.029 12.458 8.429 ;
      LAYER V1 ;
        RECT 12.338 8.166 12.438 8.266 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 11.643 10.567 12.843 10.687 ;
        RECT 12.011 8.688 12.101 10.687 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 11.643 5.787 12.843 5.907 ;
        RECT 12.011 5.787 12.101 7.721 ;
    END
  END VSS
END INVERTER

MACRO NAND
  CLASS CORE ;
  ORIGIN -11.114 -5.377 ;
  FOREIGN NAND 11.114 5.377 ;
  SIZE 1.5 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.799 7.589 11.914 7.989 ;
      LAYER M2 ;
        RECT 11.799 7.619 11.929 8.019 ;
      LAYER V1 ;
        RECT 11.808 7.756 11.908 7.856 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.099 7.589 12.214 7.989 ;
      LAYER M2 ;
        RECT 12.099 7.619 12.229 8.019 ;
      LAYER V1 ;
        RECT 12.108 7.756 12.208 7.856 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.219 8.098 12.309 9.078 ;
        RECT 11.499 8.098 12.309 8.188 ;
        RECT 11.499 7.589 11.614 7.989 ;
        RECT 11.499 6.711 11.589 9.078 ;
      LAYER M2 ;
        RECT 11.499 7.619 11.629 8.019 ;
      LAYER V1 ;
        RECT 11.509 7.756 11.609 7.856 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 11.114 10.157 12.614 10.277 ;
        RECT 11.919 8.278 12.009 10.277 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 11.114 5.377 12.614 5.497 ;
        RECT 12.219 5.377 12.309 7.311 ;
    END
  END VSS
END NAND

MACRO NOR
  CLASS CORE ;
  ORIGIN -8.994 -6.208 ;
  FOREIGN NOR 8.994 6.208 ;
  SIZE 1.8 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.279 8.438 10.394 8.832 ;
      LAYER M2 ;
        RECT 10.279 8.45 10.409 8.85 ;
      LAYER V1 ;
        RECT 10.288 8.605 10.388 8.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.679 8.438 9.794 8.832 ;
      LAYER M2 ;
        RECT 9.679 8.45 9.809 8.85 ;
      LAYER V1 ;
        RECT 9.688 8.605 9.788 8.705 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.379 8.922 9.975 9.019 ;
        RECT 9.885 7.542 9.975 9.019 ;
        RECT 9.379 8.438 9.494 8.832 ;
        RECT 9.379 8.438 9.469 9.909 ;
      LAYER M2 ;
        RECT 9.379 8.45 9.509 8.85 ;
      LAYER V1 ;
        RECT 9.389 8.605 9.489 8.705 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.994 10.988 10.794 11.108 ;
        RECT 10.399 9.109 10.489 11.108 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 8.994 6.208 10.794 6.328 ;
        RECT 10.399 6.208 10.489 8.142 ;
        RECT 9.379 6.208 9.469 8.142 ;
    END
  END VSS
END NOR

MACRO XOR
  CLASS CORE ;
  ORIGIN -12.016 -6.902 ;
  FOREIGN XOR 12.016 6.902 ;
  SIZE 3 BY 4.9 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.416 9.114 12.531 9.514 ;
      LAYER M2 ;
        RECT 12.401 9.144 12.531 9.544 ;
      LAYER V1 ;
        RECT 12.426 9.3 12.526 9.4 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.016 9.114 13.131 9.514 ;
      LAYER M2 ;
        RECT 13.001 9.144 13.131 9.544 ;
      LAYER V1 ;
        RECT 13.026 9.3 13.126 9.4 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 13.601 9.114 13.716 9.514 ;
        RECT 12.984 9.623 13.691 9.713 ;
        RECT 13.601 8.236 13.691 9.713 ;
        RECT 12.984 9.623 13.074 10.603 ;
      LAYER M2 ;
        RECT 13.601 9.144 13.731 9.544 ;
      LAYER V1 ;
        RECT 13.611 9.308 13.711 9.408 ;
    END
  END OUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT 12.016 6.902 15.016 7.022 ;
        RECT 14.616 6.902 14.706 8.836 ;
        RECT 13.928 6.902 14.018 8.836 ;
        RECT 12.38 6.902 12.47 8.836 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT 12.016 11.682 15.016 11.802 ;
        RECT 13.928 9.803 14.018 11.802 ;
    END
  END VDD
  OBS
    LAYER M1 ;
      RECT 14.616 9.623 14.706 10.603 ;
      RECT 14.316 8.234 14.406 9.715 ;
      RECT 13.808 9.623 14.706 9.713 ;
      RECT 13.808 9.126 13.92 9.713 ;
      RECT 12.38 10.984 13.54 11.074 ;
      RECT 13.45 9.803 13.54 11.074 ;
      RECT 12.38 9.803 12.47 11.074 ;
  END
END XOR

END LIBRARY
